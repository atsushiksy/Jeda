library verilog;
use verilog.vl_types.all;
entity jeda_module is
    port(
        clock           : inout  vl_logic;
        squat_rx_clk_0  : in     vl_logic;
        squat_rx_clk_1  : in     vl_logic;
        squat_rx_clk_2  : in     vl_logic;
        squat_rx_clk_3  : in     vl_logic;
        squat_rx_data_0 : out    vl_logic_vector(7 downto 0);
        squat_rx_data_1 : out    vl_logic_vector(7 downto 0);
        squat_rx_data_2 : out    vl_logic_vector(7 downto 0);
        squat_rx_data_3 : out    vl_logic_vector(7 downto 0);
        squat_rx_soc_0  : out    vl_logic;
        squat_rx_soc_1  : out    vl_logic;
        squat_rx_soc_2  : out    vl_logic;
        squat_rx_soc_3  : out    vl_logic;
        squat_rx_en_0   : in     vl_logic;
        squat_rx_en_1   : in     vl_logic;
        squat_rx_en_2   : in     vl_logic;
        squat_rx_en_3   : in     vl_logic;
        squat_rx_clav_0 : out    vl_logic;
        squat_rx_clav_1 : out    vl_logic;
        squat_rx_clav_2 : out    vl_logic;
        squat_rx_clav_3 : out    vl_logic;
        squat_tx_clk_0  : in     vl_logic;
        squat_tx_clk_1  : in     vl_logic;
        squat_tx_clk_2  : in     vl_logic;
        squat_tx_clk_3  : in     vl_logic;
        squat_tx_data_0 : in     vl_logic_vector(7 downto 0);
        squat_tx_data_1 : in     vl_logic_vector(7 downto 0);
        squat_tx_data_2 : in     vl_logic_vector(7 downto 0);
        squat_tx_data_3 : in     vl_logic_vector(7 downto 0);
        squat_tx_soc_0  : in     vl_logic;
        squat_tx_soc_1  : in     vl_logic;
        squat_tx_soc_2  : in     vl_logic;
        squat_tx_soc_3  : in     vl_logic;
        squat_tx_en_0   : in     vl_logic;
        squat_tx_en_1   : in     vl_logic;
        squat_tx_en_2   : in     vl_logic;
        squat_tx_en_3   : in     vl_logic;
        squat_tx_clav_0 : out    vl_logic;
        squat_tx_clav_1 : out    vl_logic;
        squat_tx_clav_2 : out    vl_logic;
        squat_tx_clav_3 : out    vl_logic;
        squat_busmode   : out    vl_logic;
        squat_addr      : out    vl_logic_vector(11 downto 0);
        squat_sel       : out    vl_logic;
        squat_data      : inout  vl_logic_vector(7 downto 0);
        squat_rd_ds     : out    vl_logic;
        squat_wr_rw     : out    vl_logic;
        squat_rdy_dtack : in     vl_logic;
        squat_rst       : out    vl_logic;
        squat_clk       : inout  vl_logic
    );
end jeda_module;
