library verilog;
use verilog.vl_types.all;
entity squat_test is
    generic(
        simulation_cycle: integer := 100
    );
end squat_test;
